// GENERAL DEFINITIONS
`define TRUE 1'b1
`define FALSE 1'b0

// DEFINITIONS FOR THE STATE MACHINE
`define WAITING 3'b000
`define AUTHENTICATION 3'b001
`define MENU 3'b010
`define BALANCE 3'b011
`define WITHDRAW 3'b100
`define DEPOSIT 3'b101
`define CHANGE_PIN 3'b110
`define IDLE 3'b111



// DEFINITIONS FOR THE AUTHENTICATION
`define FIND_ACCOUNT 1'b0
`define AUTHENTICATE_ACCOUNT 1'b1
`define ACCOUNT_NOT_FOUND 1'b0
`define ACCOUNT_FOUND 1'b1
`define ACCOUNT_NOT_AUTHENTICATED 1'b0
`define ACCOUNT_AUTHENTICATED 1'b1

// DEFINITIONS FOR LANGUAGE
`define ENGLISH 1'b0
`define ARABIC 1'b1